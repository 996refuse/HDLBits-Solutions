module top_module ( input a, input b, output out );
    mod_a obj(a, b, out);
endmodule
